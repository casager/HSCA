module CSAM_new (Z, X, Y);
	
	input logic [15:0] Y;
	input logic [11:0] X;
	output logic [27:0] Z;


	logic [11:0] P0;
	logic [11:0] carry1;
	logic [11:0] sum1;
	logic [11:0] P1;
	logic [11:0] carry2;
	logic [11:0] sum2;
	logic [11:0] P2;
	logic [11:0] carry3;
	logic [11:0] sum3;
	logic [11:0] P3;
	logic [11:0] carry4;
	logic [11:0] sum4;
	logic [11:0] P4;
	logic [11:0] carry5;
	logic [11:0] sum5;
	logic [11:0] P5;
	logic [11:0] carry6;
	logic [11:0] sum6;
	logic [11:0] P6;
	logic [11:0] carry7;
	logic [11:0] sum7;
	logic [11:0] P7;
	logic [11:0] carry8;
	logic [11:0] sum8;
	logic [11:0] P8;
	logic [11:0] carry9;
	logic [11:0] sum9;
	logic [11:0] P9;
	logic [11:0] carry10;
	logic [11:0] sum10;
	logic [11:0] P10;
	logic [11:0] carry11;
	logic [11:0] sum11;
	logic [11:0] P11;
	logic [11:0] carry12;
	logic [11:0] sum12;
	logic [11:0] P12;
	logic [11:0] carry13;
	logic [11:0] sum13;
	logic [11:0] P13;
	logic [11:0] carry14;
	logic [11:0] sum14;
	logic [11:0] P14;
	logic [11:0] carry15;
	logic [11:0] sum15;
	logic [11:0] P15;
	logic [11:0] carry16;
	logic [11:0] sum16;
	logic [26:0] carry17;


	// generate the partial products.
	and pp1(P0[11], X[11], Y[0]);
	and pp2(P0[10], X[10], Y[0]);
	and pp3(P0[9], X[9], Y[0]);
	and pp4(P0[8], X[8], Y[0]);
	and pp5(P0[7], X[7], Y[0]);
	and pp6(P0[6], X[6], Y[0]);
	and pp7(P0[5], X[5], Y[0]);
	and pp8(P0[4], X[4], Y[0]);
	and pp9(P0[3], X[3], Y[0]);
	and pp10(P0[2], X[2], Y[0]);
	and pp11(P0[1], X[1], Y[0]);
	and pp12(P0[0], X[0], Y[0]);
	and pp13(sum1[11], X[11], Y[1]);
	and pp14(P1[10], X[10], Y[1]);
	and pp15(P1[9], X[9], Y[1]);
	and pp16(P1[8], X[8], Y[1]);
	and pp17(P1[7], X[7], Y[1]);
	and pp18(P1[6], X[6], Y[1]);
	and pp19(P1[5], X[5], Y[1]);
	and pp20(P1[4], X[4], Y[1]);
	and pp21(P1[3], X[3], Y[1]);
	and pp22(P1[2], X[2], Y[1]);
	and pp23(P1[1], X[1], Y[1]);
	and pp24(P1[0], X[0], Y[1]);
	and pp25(sum2[11], X[11], Y[2]);
	and pp26(P2[10], X[10], Y[2]);
	and pp27(P2[9], X[9], Y[2]);
	and pp28(P2[8], X[8], Y[2]);
	and pp29(P2[7], X[7], Y[2]);
	and pp30(P2[6], X[6], Y[2]);
	and pp31(P2[5], X[5], Y[2]);
	and pp32(P2[4], X[4], Y[2]);
	and pp33(P2[3], X[3], Y[2]);
	and pp34(P2[2], X[2], Y[2]);
	and pp35(P2[1], X[1], Y[2]);
	and pp36(P2[0], X[0], Y[2]);
	and pp37(sum3[11], X[11], Y[3]);
	and pp38(P3[10], X[10], Y[3]);
	and pp39(P3[9], X[9], Y[3]);
	and pp40(P3[8], X[8], Y[3]);
	and pp41(P3[7], X[7], Y[3]);
	and pp42(P3[6], X[6], Y[3]);
	and pp43(P3[5], X[5], Y[3]);
	and pp44(P3[4], X[4], Y[3]);
	and pp45(P3[3], X[3], Y[3]);
	and pp46(P3[2], X[2], Y[3]);
	and pp47(P3[1], X[1], Y[3]);
	and pp48(P3[0], X[0], Y[3]);
	and pp49(sum4[11], X[11], Y[4]);
	and pp50(P4[10], X[10], Y[4]);
	and pp51(P4[9], X[9], Y[4]);
	and pp52(P4[8], X[8], Y[4]);
	and pp53(P4[7], X[7], Y[4]);
	and pp54(P4[6], X[6], Y[4]);
	and pp55(P4[5], X[5], Y[4]);
	and pp56(P4[4], X[4], Y[4]);
	and pp57(P4[3], X[3], Y[4]);
	and pp58(P4[2], X[2], Y[4]);
	and pp59(P4[1], X[1], Y[4]);
	and pp60(P4[0], X[0], Y[4]);
	and pp61(sum5[11], X[11], Y[5]);
	and pp62(P5[10], X[10], Y[5]);
	and pp63(P5[9], X[9], Y[5]);
	and pp64(P5[8], X[8], Y[5]);
	and pp65(P5[7], X[7], Y[5]);
	and pp66(P5[6], X[6], Y[5]);
	and pp67(P5[5], X[5], Y[5]);
	and pp68(P5[4], X[4], Y[5]);
	and pp69(P5[3], X[3], Y[5]);
	and pp70(P5[2], X[2], Y[5]);
	and pp71(P5[1], X[1], Y[5]);
	and pp72(P5[0], X[0], Y[5]);
	and pp73(sum6[11], X[11], Y[6]);
	and pp74(P6[10], X[10], Y[6]);
	and pp75(P6[9], X[9], Y[6]);
	and pp76(P6[8], X[8], Y[6]);
	and pp77(P6[7], X[7], Y[6]);
	and pp78(P6[6], X[6], Y[6]);
	and pp79(P6[5], X[5], Y[6]);
	and pp80(P6[4], X[4], Y[6]);
	and pp81(P6[3], X[3], Y[6]);
	and pp82(P6[2], X[2], Y[6]);
	and pp83(P6[1], X[1], Y[6]);
	and pp84(P6[0], X[0], Y[6]);
	and pp85(sum7[11], X[11], Y[7]);
	and pp86(P7[10], X[10], Y[7]);
	and pp87(P7[9], X[9], Y[7]);
	and pp88(P7[8], X[8], Y[7]);
	and pp89(P7[7], X[7], Y[7]);
	and pp90(P7[6], X[6], Y[7]);
	and pp91(P7[5], X[5], Y[7]);
	and pp92(P7[4], X[4], Y[7]);
	and pp93(P7[3], X[3], Y[7]);
	and pp94(P7[2], X[2], Y[7]);
	and pp95(P7[1], X[1], Y[7]);
	and pp96(P7[0], X[0], Y[7]);
	and pp97(sum8[11], X[11], Y[8]);
	and pp98(P8[10], X[10], Y[8]);
	and pp99(P8[9], X[9], Y[8]);
	and pp100(P8[8], X[8], Y[8]);
	and pp101(P8[7], X[7], Y[8]);
	and pp102(P8[6], X[6], Y[8]);
	and pp103(P8[5], X[5], Y[8]);
	and pp104(P8[4], X[4], Y[8]);
	and pp105(P8[3], X[3], Y[8]);
	and pp106(P8[2], X[2], Y[8]);
	and pp107(P8[1], X[1], Y[8]);
	and pp108(P8[0], X[0], Y[8]);
	and pp109(sum9[11], X[11], Y[9]);
	and pp110(P9[10], X[10], Y[9]);
	and pp111(P9[9], X[9], Y[9]);
	and pp112(P9[8], X[8], Y[9]);
	and pp113(P9[7], X[7], Y[9]);
	and pp114(P9[6], X[6], Y[9]);
	and pp115(P9[5], X[5], Y[9]);
	and pp116(P9[4], X[4], Y[9]);
	and pp117(P9[3], X[3], Y[9]);
	and pp118(P9[2], X[2], Y[9]);
	and pp119(P9[1], X[1], Y[9]);
	and pp120(P9[0], X[0], Y[9]);
	and pp121(sum10[11], X[11], Y[10]);
	and pp122(P10[10], X[10], Y[10]);
	and pp123(P10[9], X[9], Y[10]);
	and pp124(P10[8], X[8], Y[10]);
	and pp125(P10[7], X[7], Y[10]);
	and pp126(P10[6], X[6], Y[10]);
	and pp127(P10[5], X[5], Y[10]);
	and pp128(P10[4], X[4], Y[10]);
	and pp129(P10[3], X[3], Y[10]);
	and pp130(P10[2], X[2], Y[10]);
	and pp131(P10[1], X[1], Y[10]);
	and pp132(P10[0], X[0], Y[10]);
	and pp133(sum11[11], X[11], Y[11]);
	and pp134(P11[10], X[10], Y[11]);
	and pp135(P11[9], X[9], Y[11]);
	and pp136(P11[8], X[8], Y[11]);
	and pp137(P11[7], X[7], Y[11]);
	and pp138(P11[6], X[6], Y[11]);
	and pp139(P11[5], X[5], Y[11]);
	and pp140(P11[4], X[4], Y[11]);
	and pp141(P11[3], X[3], Y[11]);
	and pp142(P11[2], X[2], Y[11]);
	and pp143(P11[1], X[1], Y[11]);
	and pp144(P11[0], X[0], Y[11]);
	and pp145(sum12[11], X[11], Y[12]);
	and pp146(P12[10], X[10], Y[12]);
	and pp147(P12[9], X[9], Y[12]);
	and pp148(P12[8], X[8], Y[12]);
	and pp149(P12[7], X[7], Y[12]);
	and pp150(P12[6], X[6], Y[12]);
	and pp151(P12[5], X[5], Y[12]);
	and pp152(P12[4], X[4], Y[12]);
	and pp153(P12[3], X[3], Y[12]);
	and pp154(P12[2], X[2], Y[12]);
	and pp155(P12[1], X[1], Y[12]);
	and pp156(P12[0], X[0], Y[12]);
	and pp157(sum13[11], X[11], Y[13]);
	and pp158(P13[10], X[10], Y[13]);
	and pp159(P13[9], X[9], Y[13]);
	and pp160(P13[8], X[8], Y[13]);
	and pp161(P13[7], X[7], Y[13]);
	and pp162(P13[6], X[6], Y[13]);
	and pp163(P13[5], X[5], Y[13]);
	and pp164(P13[4], X[4], Y[13]);
	and pp165(P13[3], X[3], Y[13]);
	and pp166(P13[2], X[2], Y[13]);
	and pp167(P13[1], X[1], Y[13]);
	and pp168(P13[0], X[0], Y[13]);
	and pp169(sum14[11], X[11], Y[14]);
	and pp170(P14[10], X[10], Y[14]);
	and pp171(P14[9], X[9], Y[14]);
	and pp172(P14[8], X[8], Y[14]);
	and pp173(P14[7], X[7], Y[14]);
	and pp174(P14[6], X[6], Y[14]);
	and pp175(P14[5], X[5], Y[14]);
	and pp176(P14[4], X[4], Y[14]);
	and pp177(P14[3], X[3], Y[14]);
	and pp178(P14[2], X[2], Y[14]);
	and pp179(P14[1], X[1], Y[14]);
	and pp180(P14[0], X[0], Y[14]);
	and pp181(sum15[11], X[11], Y[15]);
	and pp182(P15[10], X[10], Y[15]);
	and pp183(P15[9], X[9], Y[15]);
	and pp184(P15[8], X[8], Y[15]);
	and pp185(P15[7], X[7], Y[15]);
	and pp186(P15[6], X[6], Y[15]);
	and pp187(P15[5], X[5], Y[15]);
	and pp188(P15[4], X[4], Y[15]);
	and pp189(P15[3], X[3], Y[15]);
	and pp190(P15[2], X[2], Y[15]);
	and pp191(P15[1], X[1], Y[15]);
	and pp192(P15[0], X[0], Y[15]);

	// Array Reduction
	half_adder  HA1(carry1[10],sum1[10],P1[10],P0[11]);
	half_adder  HA2(carry1[9],sum1[9],P1[9],P0[10]);
	half_adder  HA3(carry1[8],sum1[8],P1[8],P0[9]);
	half_adder  HA4(carry1[7],sum1[7],P1[7],P0[8]);
	half_adder  HA5(carry1[6],sum1[6],P1[6],P0[7]);
	half_adder  HA6(carry1[5],sum1[5],P1[5],P0[6]);
	half_adder  HA7(carry1[4],sum1[4],P1[4],P0[5]);
	half_adder  HA8(carry1[3],sum1[3],P1[3],P0[4]);
	half_adder  HA9(carry1[2],sum1[2],P1[2],P0[3]);
	half_adder  HA10(carry1[1],sum1[1],P1[1],P0[2]);
	half_adder  HA11(carry1[0],sum1[0],P1[0],P0[1]);
	full_adder  FA1(carry2[10],sum2[10],P2[10],sum1[11],carry1[10]);
	full_adder  FA2(carry2[9],sum2[9],P2[9],sum1[10],carry1[9]);
	full_adder  FA3(carry2[8],sum2[8],P2[8],sum1[9],carry1[8]);
	full_adder  FA4(carry2[7],sum2[7],P2[7],sum1[8],carry1[7]);
	full_adder  FA5(carry2[6],sum2[6],P2[6],sum1[7],carry1[6]);
	full_adder  FA6(carry2[5],sum2[5],P2[5],sum1[6],carry1[5]);
	full_adder  FA7(carry2[4],sum2[4],P2[4],sum1[5],carry1[4]);
	full_adder  FA8(carry2[3],sum2[3],P2[3],sum1[4],carry1[3]);
	full_adder  FA9(carry2[2],sum2[2],P2[2],sum1[3],carry1[2]);
	full_adder  FA10(carry2[1],sum2[1],P2[1],sum1[2],carry1[1]);
	full_adder  FA11(carry2[0],sum2[0],P2[0],sum1[1],carry1[0]);
	full_adder  FA12(carry3[10],sum3[10],P3[10],sum2[11],carry2[10]);
	full_adder  FA13(carry3[9],sum3[9],P3[9],sum2[10],carry2[9]);
	full_adder  FA14(carry3[8],sum3[8],P3[8],sum2[9],carry2[8]);
	full_adder  FA15(carry3[7],sum3[7],P3[7],sum2[8],carry2[7]);
	full_adder  FA16(carry3[6],sum3[6],P3[6],sum2[7],carry2[6]);
	full_adder  FA17(carry3[5],sum3[5],P3[5],sum2[6],carry2[5]);
	full_adder  FA18(carry3[4],sum3[4],P3[4],sum2[5],carry2[4]);
	full_adder  FA19(carry3[3],sum3[3],P3[3],sum2[4],carry2[3]);
	full_adder  FA20(carry3[2],sum3[2],P3[2],sum2[3],carry2[2]);
	full_adder  FA21(carry3[1],sum3[1],P3[1],sum2[2],carry2[1]);
	full_adder  FA22(carry3[0],sum3[0],P3[0],sum2[1],carry2[0]);
	full_adder  FA23(carry4[10],sum4[10],P4[10],sum3[11],carry3[10]);
	full_adder  FA24(carry4[9],sum4[9],P4[9],sum3[10],carry3[9]);
	full_adder  FA25(carry4[8],sum4[8],P4[8],sum3[9],carry3[8]);
	full_adder  FA26(carry4[7],sum4[7],P4[7],sum3[8],carry3[7]);
	full_adder  FA27(carry4[6],sum4[6],P4[6],sum3[7],carry3[6]);
	full_adder  FA28(carry4[5],sum4[5],P4[5],sum3[6],carry3[5]);
	full_adder  FA29(carry4[4],sum4[4],P4[4],sum3[5],carry3[4]);
	full_adder  FA30(carry4[3],sum4[3],P4[3],sum3[4],carry3[3]);
	full_adder  FA31(carry4[2],sum4[2],P4[2],sum3[3],carry3[2]);
	full_adder  FA32(carry4[1],sum4[1],P4[1],sum3[2],carry3[1]);
	full_adder  FA33(carry4[0],sum4[0],P4[0],sum3[1],carry3[0]);
	full_adder  FA34(carry5[10],sum5[10],P5[10],sum4[11],carry4[10]);
	full_adder  FA35(carry5[9],sum5[9],P5[9],sum4[10],carry4[9]);
	full_adder  FA36(carry5[8],sum5[8],P5[8],sum4[9],carry4[8]);
	full_adder  FA37(carry5[7],sum5[7],P5[7],sum4[8],carry4[7]);
	full_adder  FA38(carry5[6],sum5[6],P5[6],sum4[7],carry4[6]);
	full_adder  FA39(carry5[5],sum5[5],P5[5],sum4[6],carry4[5]);
	full_adder  FA40(carry5[4],sum5[4],P5[4],sum4[5],carry4[4]);
	full_adder  FA41(carry5[3],sum5[3],P5[3],sum4[4],carry4[3]);
	full_adder  FA42(carry5[2],sum5[2],P5[2],sum4[3],carry4[2]);
	full_adder  FA43(carry5[1],sum5[1],P5[1],sum4[2],carry4[1]);
	full_adder  FA44(carry5[0],sum5[0],P5[0],sum4[1],carry4[0]);
	full_adder  FA45(carry6[10],sum6[10],P6[10],sum5[11],carry5[10]);
	full_adder  FA46(carry6[9],sum6[9],P6[9],sum5[10],carry5[9]);
	full_adder  FA47(carry6[8],sum6[8],P6[8],sum5[9],carry5[8]);
	full_adder  FA48(carry6[7],sum6[7],P6[7],sum5[8],carry5[7]);
	full_adder  FA49(carry6[6],sum6[6],P6[6],sum5[7],carry5[6]);
	full_adder  FA50(carry6[5],sum6[5],P6[5],sum5[6],carry5[5]);
	full_adder  FA51(carry6[4],sum6[4],P6[4],sum5[5],carry5[4]);
	full_adder  FA52(carry6[3],sum6[3],P6[3],sum5[4],carry5[3]);
	full_adder  FA53(carry6[2],sum6[2],P6[2],sum5[3],carry5[2]);
	full_adder  FA54(carry6[1],sum6[1],P6[1],sum5[2],carry5[1]);
	full_adder  FA55(carry6[0],sum6[0],P6[0],sum5[1],carry5[0]);
	full_adder  FA56(carry7[10],sum7[10],P7[10],sum6[11],carry6[10]);
	full_adder  FA57(carry7[9],sum7[9],P7[9],sum6[10],carry6[9]);
	full_adder  FA58(carry7[8],sum7[8],P7[8],sum6[9],carry6[8]);
	full_adder  FA59(carry7[7],sum7[7],P7[7],sum6[8],carry6[7]);
	full_adder  FA60(carry7[6],sum7[6],P7[6],sum6[7],carry6[6]);
	full_adder  FA61(carry7[5],sum7[5],P7[5],sum6[6],carry6[5]);
	full_adder  FA62(carry7[4],sum7[4],P7[4],sum6[5],carry6[4]);
	full_adder  FA63(carry7[3],sum7[3],P7[3],sum6[4],carry6[3]);
	full_adder  FA64(carry7[2],sum7[2],P7[2],sum6[3],carry6[2]);
	full_adder  FA65(carry7[1],sum7[1],P7[1],sum6[2],carry6[1]);
	full_adder  FA66(carry7[0],sum7[0],P7[0],sum6[1],carry6[0]);
	full_adder  FA67(carry8[10],sum8[10],P8[10],sum7[11],carry7[10]);
	full_adder  FA68(carry8[9],sum8[9],P8[9],sum7[10],carry7[9]);
	full_adder  FA69(carry8[8],sum8[8],P8[8],sum7[9],carry7[8]);
	full_adder  FA70(carry8[7],sum8[7],P8[7],sum7[8],carry7[7]);
	full_adder  FA71(carry8[6],sum8[6],P8[6],sum7[7],carry7[6]);
	full_adder  FA72(carry8[5],sum8[5],P8[5],sum7[6],carry7[5]);
	full_adder  FA73(carry8[4],sum8[4],P8[4],sum7[5],carry7[4]);
	full_adder  FA74(carry8[3],sum8[3],P8[3],sum7[4],carry7[3]);
	full_adder  FA75(carry8[2],sum8[2],P8[2],sum7[3],carry7[2]);
	full_adder  FA76(carry8[1],sum8[1],P8[1],sum7[2],carry7[1]);
	full_adder  FA77(carry8[0],sum8[0],P8[0],sum7[1],carry7[0]);
	full_adder  FA78(carry9[10],sum9[10],P9[10],sum8[11],carry8[10]);
	full_adder  FA79(carry9[9],sum9[9],P9[9],sum8[10],carry8[9]);
	full_adder  FA80(carry9[8],sum9[8],P9[8],sum8[9],carry8[8]);
	full_adder  FA81(carry9[7],sum9[7],P9[7],sum8[8],carry8[7]);
	full_adder  FA82(carry9[6],sum9[6],P9[6],sum8[7],carry8[6]);
	full_adder  FA83(carry9[5],sum9[5],P9[5],sum8[6],carry8[5]);
	full_adder  FA84(carry9[4],sum9[4],P9[4],sum8[5],carry8[4]);
	full_adder  FA85(carry9[3],sum9[3],P9[3],sum8[4],carry8[3]);
	full_adder  FA86(carry9[2],sum9[2],P9[2],sum8[3],carry8[2]);
	full_adder  FA87(carry9[1],sum9[1],P9[1],sum8[2],carry8[1]);
	full_adder  FA88(carry9[0],sum9[0],P9[0],sum8[1],carry8[0]);
	full_adder  FA89(carry10[10],sum10[10],P10[10],sum9[11],carry9[10]);
	full_adder  FA90(carry10[9],sum10[9],P10[9],sum9[10],carry9[9]);
	full_adder  FA91(carry10[8],sum10[8],P10[8],sum9[9],carry9[8]);
	full_adder  FA92(carry10[7],sum10[7],P10[7],sum9[8],carry9[7]);
	full_adder  FA93(carry10[6],sum10[6],P10[6],sum9[7],carry9[6]);
	full_adder  FA94(carry10[5],sum10[5],P10[5],sum9[6],carry9[5]);
	full_adder  FA95(carry10[4],sum10[4],P10[4],sum9[5],carry9[4]);
	full_adder  FA96(carry10[3],sum10[3],P10[3],sum9[4],carry9[3]);
	full_adder  FA97(carry10[2],sum10[2],P10[2],sum9[3],carry9[2]);
	full_adder  FA98(carry10[1],sum10[1],P10[1],sum9[2],carry9[1]);
	full_adder  FA99(carry10[0],sum10[0],P10[0],sum9[1],carry9[0]);
	full_adder  FA100(carry11[10],sum11[10],P11[10],sum10[11],carry10[10]);
	full_adder  FA101(carry11[9],sum11[9],P11[9],sum10[10],carry10[9]);
	full_adder  FA102(carry11[8],sum11[8],P11[8],sum10[9],carry10[8]);
	full_adder  FA103(carry11[7],sum11[7],P11[7],sum10[8],carry10[7]);
	full_adder  FA104(carry11[6],sum11[6],P11[6],sum10[7],carry10[6]);
	full_adder  FA105(carry11[5],sum11[5],P11[5],sum10[6],carry10[5]);
	full_adder  FA106(carry11[4],sum11[4],P11[4],sum10[5],carry10[4]);
	full_adder  FA107(carry11[3],sum11[3],P11[3],sum10[4],carry10[3]);
	full_adder  FA108(carry11[2],sum11[2],P11[2],sum10[3],carry10[2]);
	full_adder  FA109(carry11[1],sum11[1],P11[1],sum10[2],carry10[1]);
	full_adder  FA110(carry11[0],sum11[0],P11[0],sum10[1],carry10[0]);
	full_adder  FA111(carry12[10],sum12[10],P12[10],sum11[11],carry11[10]);
	full_adder  FA112(carry12[9],sum12[9],P12[9],sum11[10],carry11[9]);
	full_adder  FA113(carry12[8],sum12[8],P12[8],sum11[9],carry11[8]);
	full_adder  FA114(carry12[7],sum12[7],P12[7],sum11[8],carry11[7]);
	full_adder  FA115(carry12[6],sum12[6],P12[6],sum11[7],carry11[6]);
	full_adder  FA116(carry12[5],sum12[5],P12[5],sum11[6],carry11[5]);
	full_adder  FA117(carry12[4],sum12[4],P12[4],sum11[5],carry11[4]);
	full_adder  FA118(carry12[3],sum12[3],P12[3],sum11[4],carry11[3]);
	full_adder  FA119(carry12[2],sum12[2],P12[2],sum11[3],carry11[2]);
	full_adder  FA120(carry12[1],sum12[1],P12[1],sum11[2],carry11[1]);
	full_adder  FA121(carry12[0],sum12[0],P12[0],sum11[1],carry11[0]);
	full_adder  FA122(carry13[10],sum13[10],P13[10],sum12[11],carry12[10]);
	full_adder  FA123(carry13[9],sum13[9],P13[9],sum12[10],carry12[9]);
	full_adder  FA124(carry13[8],sum13[8],P13[8],sum12[9],carry12[8]);
	full_adder  FA125(carry13[7],sum13[7],P13[7],sum12[8],carry12[7]);
	full_adder  FA126(carry13[6],sum13[6],P13[6],sum12[7],carry12[6]);
	full_adder  FA127(carry13[5],sum13[5],P13[5],sum12[6],carry12[5]);
	full_adder  FA128(carry13[4],sum13[4],P13[4],sum12[5],carry12[4]);
	full_adder  FA129(carry13[3],sum13[3],P13[3],sum12[4],carry12[3]);
	full_adder  FA130(carry13[2],sum13[2],P13[2],sum12[3],carry12[2]);
	full_adder  FA131(carry13[1],sum13[1],P13[1],sum12[2],carry12[1]);
	full_adder  FA132(carry13[0],sum13[0],P13[0],sum12[1],carry12[0]);
	full_adder  FA133(carry14[10],sum14[10],P14[10],sum13[11],carry13[10]);
	full_adder  FA134(carry14[9],sum14[9],P14[9],sum13[10],carry13[9]);
	full_adder  FA135(carry14[8],sum14[8],P14[8],sum13[9],carry13[8]);
	full_adder  FA136(carry14[7],sum14[7],P14[7],sum13[8],carry13[7]);
	full_adder  FA137(carry14[6],sum14[6],P14[6],sum13[7],carry13[6]);
	full_adder  FA138(carry14[5],sum14[5],P14[5],sum13[6],carry13[5]);
	full_adder  FA139(carry14[4],sum14[4],P14[4],sum13[5],carry13[4]);
	full_adder  FA140(carry14[3],sum14[3],P14[3],sum13[4],carry13[3]);
	full_adder  FA141(carry14[2],sum14[2],P14[2],sum13[3],carry13[2]);
	full_adder  FA142(carry14[1],sum14[1],P14[1],sum13[2],carry13[1]);
	full_adder  FA143(carry14[0],sum14[0],P14[0],sum13[1],carry13[0]);
	full_adder  FA144(carry15[10],sum15[10],P15[10],sum14[11],carry14[10]);
	full_adder  FA145(carry15[9],sum15[9],P15[9],sum14[10],carry14[9]);
	full_adder  FA146(carry15[8],sum15[8],P15[8],sum14[9],carry14[8]);
	full_adder  FA147(carry15[7],sum15[7],P15[7],sum14[8],carry14[7]);
	full_adder  FA148(carry15[6],sum15[6],P15[6],sum14[7],carry14[6]);
	full_adder  FA149(carry15[5],sum15[5],P15[5],sum14[6],carry14[5]);
	full_adder  FA150(carry15[4],sum15[4],P15[4],sum14[5],carry14[4]);
	full_adder  FA151(carry15[3],sum15[3],P15[3],sum14[4],carry14[3]);
	full_adder  FA152(carry15[2],sum15[2],P15[2],sum14[3],carry14[2]);
	full_adder  FA153(carry15[1],sum15[1],P15[1],sum14[2],carry14[1]);
	full_adder  FA154(carry15[0],sum15[0],P15[0],sum14[1],carry14[0]);

	// Generate lower product bits YBITS 
	buf b1(Z[0], P0[0]);
	assign Z[1] = sum1[0];
	assign Z[2] = sum2[0];
	assign Z[3] = sum3[0];
	assign Z[4] = sum4[0];
	assign Z[5] = sum5[0];
	assign Z[6] = sum6[0];
	assign Z[7] = sum7[0];
	assign Z[8] = sum8[0];
	assign Z[9] = sum9[0];
	assign Z[10] = sum10[0];
	assign Z[11] = sum11[0];
	assign Z[12] = sum12[0];
	assign Z[13] = sum13[0];
	assign Z[14] = sum14[0];
	assign Z[15] = sum15[0];

	// Final Carry Propagate Addition
	half_adder CPA1(carry16[0],Z[16],carry15[0],sum15[1]);
	full_adder CPA2(carry16[1],Z[17],carry15[1],carry16[0],sum15[2]);
	full_adder CPA3(carry16[2],Z[18],carry15[2],carry16[1],sum15[3]);
	full_adder CPA4(carry16[3],Z[19],carry15[3],carry16[2],sum15[4]);
	full_adder CPA5(carry16[4],Z[20],carry15[4],carry16[3],sum15[5]);
	full_adder CPA6(carry16[5],Z[21],carry15[5],carry16[4],sum15[6]);
	full_adder CPA7(carry16[6],Z[22],carry15[6],carry16[5],sum15[7]);
	full_adder CPA8(carry16[7],Z[23],carry15[7],carry16[6],sum15[8]);
	full_adder CPA9(carry16[8],Z[24],carry15[8],carry16[7],sum15[9]);
	full_adder CPA10(carry16[9],Z[25],carry15[9],carry16[8],sum15[10]);
	full_adder CPA11(Z[27],Z[26],carry15[10],carry16[9],sum15[11]);

endmodule
